magic
tech sky130A
magscale 1 2
timestamp 1672556029
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2048 178848 117552
<< metal2 >>
rect 11334 119200 11390 120000
rect 33782 119200 33838 120000
rect 56230 119200 56286 120000
rect 78678 119200 78734 120000
rect 101126 119200 101182 120000
rect 123574 119200 123630 120000
rect 146022 119200 146078 120000
rect 168470 119200 168526 120000
rect 5446 0 5502 800
rect 15382 0 15438 800
rect 25318 0 25374 800
rect 35254 0 35310 800
rect 45190 0 45246 800
rect 55126 0 55182 800
rect 65062 0 65118 800
rect 74998 0 75054 800
rect 84934 0 84990 800
rect 94870 0 94926 800
rect 104806 0 104862 800
rect 114742 0 114798 800
rect 124678 0 124734 800
rect 134614 0 134670 800
rect 144550 0 144606 800
rect 154486 0 154542 800
rect 164422 0 164478 800
rect 174358 0 174414 800
<< obsm2 >>
rect 4214 119144 11278 119354
rect 11446 119144 33726 119354
rect 33894 119144 56174 119354
rect 56342 119144 78622 119354
rect 78790 119144 101070 119354
rect 101238 119144 123518 119354
rect 123686 119144 145966 119354
rect 146134 119144 168414 119354
rect 168582 119144 174412 119354
rect 4214 856 174412 119144
rect 4214 734 5390 856
rect 5558 734 15326 856
rect 15494 734 25262 856
rect 25430 734 35198 856
rect 35366 734 45134 856
rect 45302 734 55070 856
rect 55238 734 65006 856
rect 65174 734 74942 856
rect 75110 734 84878 856
rect 85046 734 94814 856
rect 94982 734 104750 856
rect 104918 734 114686 856
rect 114854 734 124622 856
rect 124790 734 134558 856
rect 134726 734 144494 856
rect 144662 734 154430 856
rect 154598 734 164366 856
rect 164534 734 174302 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 25318 0 25374 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 A[1]
port 2 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 A[2]
port 3 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 A[3]
port 4 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 A[4]
port 5 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 A[5]
port 6 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 A[6]
port 7 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 A[7]
port 8 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 B[0]
port 9 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 B[1]
port 10 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 B[2]
port 11 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 B[3]
port 12 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 B[4]
port 13 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 B[5]
port 14 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 B[6]
port 15 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 B[7]
port 16 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 clock
port 17 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 reset
port 18 nsew signal input
rlabel metal2 s 11334 119200 11390 120000 6 sum[0]
port 19 nsew signal output
rlabel metal2 s 33782 119200 33838 120000 6 sum[1]
port 20 nsew signal output
rlabel metal2 s 56230 119200 56286 120000 6 sum[2]
port 21 nsew signal output
rlabel metal2 s 78678 119200 78734 120000 6 sum[3]
port 22 nsew signal output
rlabel metal2 s 101126 119200 101182 120000 6 sum[4]
port 23 nsew signal output
rlabel metal2 s 123574 119200 123630 120000 6 sum[5]
port 24 nsew signal output
rlabel metal2 s 146022 119200 146078 120000 6 sum[6]
port 25 nsew signal output
rlabel metal2 s 168470 119200 168526 120000 6 sum[7]
port 26 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5863058
string GDS_FILE /home/rakshith/Numerical_method_bisection/openlane/user_proj_example/runs/23_01_01_12_21/results/signoff/user_proj_example.magic.gds
string GDS_START 219076
<< end >>

